��  CCircuit��  CSerializeHack           ��  CPart              ��� 
 CCapacitor��  CValue  ����    10nF(    :�0�yE>      �?nF �� 	 CTerminal  ����         ������
@          �  ����                            ����        ��      �t(gL�a>��  CECapacitor
�  � ��    470�F(    !�J�>?      �?�F �  (�)�         C�q�ut?      �;  �  (�)�                      ��    �4�        ��      !������>�� 
 CVoltmeter��  CMeter  ���     0.00(    �   �!�                �          �   �!�                            �,�        ��      ��  CEarth�  ()%                 ���fo?    $3,         ��      ��  C555�  �H�]               @N贁Nk?  �  �H�]               @          �  h`}a        C�q�ut?��'^@?  �  hp}q        C�q�ut?          �  h�}�              @          �  ����                ���fo�  �  ����        ������
@      �;  �  �p�q               �            |\��         ��   (   �� 	 CResistor
�  #'    10k          ��@      �?k  �  ( )               @��'^@?  �  (,)A        C�q�ut?��'^@�    $,,     *    ��      ��  CSPST��  CToggle  � � 0     -   �  � ,� A              @          �  �  �        	       @            � � ,    0     ��    �� 	 CVoltRail
�  [ � �     5V(          @      �? V �  �  �               @���fo�    � � �      5    ����                   ���  CWire�� 
 CCrossOver  &|,�        (p)�       7�  (`)q       7�  (piq      7�  (�)       7�9�  &|,�        � �i�      7�  �  )      7�  (`ia      7�  (@)a       7�  � @� �       7�  �p!q      7�   p!�       7�  ���       7�  �!      7�   �!       7�  ��      7�  ����       7�  ����      7�  ���       7�  (�      7�  � �      7�  ( �      7�  � �I       7�  � �I                     ���  CProbe  )�8�      8        S�  �a�p       D                                     K    F  8    =  E    H  M   Q    P   ! A ! " < " # > # $ $ L % % J & & D * @ * + + B 0 0 C 1 @ 1 5 5 1 8 ? ;  B < 8 "   > : C # 5 O ; ! + A 0 > & E D   I F H  G L G % K J  $ M = I O Q * P N   N            �$s�        @     +        @            @    "V  (      �               
         @      �? V       �      �? V         
         $@      �? V               �? V                 @      �? s 